// 4-bit encoding for each lo_discount value
// 512-way parallelism

module discount_sumv2
   (
    input  logic clk,
    
    input  logic reset,
    input  logic en,
              
    input  logic [511:0] discount_cl [3:0], // lo_discount block    
    input  logic [511:0] bit_map, // d_year scan result
        
    output logic [511:0] agg_result [3:0], // pre-reduce
    output logic processing_done
    );
		
	always_ff @(posedge clk)
	begin		
		if (reset)	
		begin				
			processing_done <= 1'b0;		
		end
		else if (en)
		begin
			agg_result[0] <= discount_cl[0] * bit_map[0];
			agg_result[1] <= discount_cl[1] * bit_map[1];
			agg_result[2] <= discount_cl[2] * bit_map[2];
			agg_result[3] <= discount_cl[3] * bit_map[3];
			agg_result[4] <= discount_cl[4] * bit_map[4];
			agg_result[5] <= discount_cl[5] * bit_map[5];
			agg_result[6] <= discount_cl[6] * bit_map[6];
			agg_result[7] <= discount_cl[7] * bit_map[7];
			agg_result[8] <= discount_cl[8] * bit_map[8];
			agg_result[9] <= discount_cl[9] * bit_map[9];
			agg_result[10] <= discount_cl[10] * bit_map[10];
			agg_result[11] <= discount_cl[11] * bit_map[11];
			agg_result[12] <= discount_cl[12] * bit_map[12];
			agg_result[13] <= discount_cl[13] * bit_map[13];
			agg_result[14] <= discount_cl[14] * bit_map[14];
			agg_result[15] <= discount_cl[15] * bit_map[15];
			agg_result[16] <= discount_cl[16] * bit_map[16];
			agg_result[17] <= discount_cl[17] * bit_map[17];
			agg_result[18] <= discount_cl[18] * bit_map[18];
			agg_result[19] <= discount_cl[19] * bit_map[19];
			agg_result[20] <= discount_cl[20] * bit_map[20];
			agg_result[21] <= discount_cl[21] * bit_map[21];
			agg_result[22] <= discount_cl[22] * bit_map[22];
			agg_result[23] <= discount_cl[23] * bit_map[23];
			agg_result[24] <= discount_cl[24] * bit_map[24];
			agg_result[25] <= discount_cl[25] * bit_map[25];
			agg_result[26] <= discount_cl[26] * bit_map[26];
			agg_result[27] <= discount_cl[27] * bit_map[27];
			agg_result[28] <= discount_cl[28] * bit_map[28];
			agg_result[29] <= discount_cl[29] * bit_map[29];
			agg_result[30] <= discount_cl[30] * bit_map[30];
			agg_result[31] <= discount_cl[31] * bit_map[31];
			agg_result[32] <= discount_cl[32] * bit_map[32];
			agg_result[33] <= discount_cl[33] * bit_map[33];
			agg_result[34] <= discount_cl[34] * bit_map[34];
			agg_result[35] <= discount_cl[35] * bit_map[35];
			agg_result[36] <= discount_cl[36] * bit_map[36];
			agg_result[37] <= discount_cl[37] * bit_map[37];
			agg_result[38] <= discount_cl[38] * bit_map[38];
			agg_result[39] <= discount_cl[39] * bit_map[39];
			agg_result[40] <= discount_cl[40] * bit_map[40];
			agg_result[41] <= discount_cl[41] * bit_map[41];
			agg_result[42] <= discount_cl[42] * bit_map[42];
			agg_result[43] <= discount_cl[43] * bit_map[43];
			agg_result[44] <= discount_cl[44] * bit_map[44];
			agg_result[45] <= discount_cl[45] * bit_map[45];
			agg_result[46] <= discount_cl[46] * bit_map[46];
			agg_result[47] <= discount_cl[47] * bit_map[47];
			agg_result[48] <= discount_cl[48] * bit_map[48];
			agg_result[49] <= discount_cl[49] * bit_map[49];
			agg_result[50] <= discount_cl[50] * bit_map[50];
			agg_result[51] <= discount_cl[51] * bit_map[51];
			agg_result[52] <= discount_cl[52] * bit_map[52];
			agg_result[53] <= discount_cl[53] * bit_map[53];
			agg_result[54] <= discount_cl[54] * bit_map[54];
			agg_result[55] <= discount_cl[55] * bit_map[55];
			agg_result[56] <= discount_cl[56] * bit_map[56];
			agg_result[57] <= discount_cl[57] * bit_map[57];
			agg_result[58] <= discount_cl[58] * bit_map[58];
			agg_result[59] <= discount_cl[59] * bit_map[59];
			agg_result[60] <= discount_cl[60] * bit_map[60];
			agg_result[61] <= discount_cl[61] * bit_map[61];
			agg_result[62] <= discount_cl[62] * bit_map[62];
			agg_result[63] <= discount_cl[63] * bit_map[63];
			agg_result[64] <= discount_cl[64] * bit_map[64];
			agg_result[65] <= discount_cl[65] * bit_map[65];
			agg_result[66] <= discount_cl[66] * bit_map[66];
			agg_result[67] <= discount_cl[67] * bit_map[67];
			agg_result[68] <= discount_cl[68] * bit_map[68];
			agg_result[69] <= discount_cl[69] * bit_map[69];
			agg_result[70] <= discount_cl[70] * bit_map[70];
			agg_result[71] <= discount_cl[71] * bit_map[71];
			agg_result[72] <= discount_cl[72] * bit_map[72];
			agg_result[73] <= discount_cl[73] * bit_map[73];
			agg_result[74] <= discount_cl[74] * bit_map[74];
			agg_result[75] <= discount_cl[75] * bit_map[75];
			agg_result[76] <= discount_cl[76] * bit_map[76];
			agg_result[77] <= discount_cl[77] * bit_map[77];
			agg_result[78] <= discount_cl[78] * bit_map[78];
			agg_result[79] <= discount_cl[79] * bit_map[79];
			agg_result[80] <= discount_cl[80] * bit_map[80];
			agg_result[81] <= discount_cl[81] * bit_map[81];
			agg_result[82] <= discount_cl[82] * bit_map[82];
			agg_result[83] <= discount_cl[83] * bit_map[83];
			agg_result[84] <= discount_cl[84] * bit_map[84];
			agg_result[85] <= discount_cl[85] * bit_map[85];
			agg_result[86] <= discount_cl[86] * bit_map[86];
			agg_result[87] <= discount_cl[87] * bit_map[87];
			agg_result[88] <= discount_cl[88] * bit_map[88];
			agg_result[89] <= discount_cl[89] * bit_map[89];
			agg_result[90] <= discount_cl[90] * bit_map[90];
			agg_result[91] <= discount_cl[91] * bit_map[91];
			agg_result[92] <= discount_cl[92] * bit_map[92];
			agg_result[93] <= discount_cl[93] * bit_map[93];
			agg_result[94] <= discount_cl[94] * bit_map[94];
			agg_result[95] <= discount_cl[95] * bit_map[95];
			agg_result[96] <= discount_cl[96] * bit_map[96];
			agg_result[97] <= discount_cl[97] * bit_map[97];
			agg_result[98] <= discount_cl[98] * bit_map[98];
			agg_result[99] <= discount_cl[99] * bit_map[99];
			agg_result[100] <= discount_cl[100] * bit_map[100];
			agg_result[101] <= discount_cl[101] * bit_map[101];
			agg_result[102] <= discount_cl[102] * bit_map[102];
			agg_result[103] <= discount_cl[103] * bit_map[103];
			agg_result[104] <= discount_cl[104] * bit_map[104];
			agg_result[105] <= discount_cl[105] * bit_map[105];
			agg_result[106] <= discount_cl[106] * bit_map[106];
			agg_result[107] <= discount_cl[107] * bit_map[107];
			agg_result[108] <= discount_cl[108] * bit_map[108];
			agg_result[109] <= discount_cl[109] * bit_map[109];
			agg_result[110] <= discount_cl[110] * bit_map[110];
			agg_result[111] <= discount_cl[111] * bit_map[111];
			agg_result[112] <= discount_cl[112] * bit_map[112];
			agg_result[113] <= discount_cl[113] * bit_map[113];
			agg_result[114] <= discount_cl[114] * bit_map[114];
			agg_result[115] <= discount_cl[115] * bit_map[115];
			agg_result[116] <= discount_cl[116] * bit_map[116];
			agg_result[117] <= discount_cl[117] * bit_map[117];
			agg_result[118] <= discount_cl[118] * bit_map[118];
			agg_result[119] <= discount_cl[119] * bit_map[119];
			agg_result[120] <= discount_cl[120] * bit_map[120];
			agg_result[121] <= discount_cl[121] * bit_map[121];
			agg_result[122] <= discount_cl[122] * bit_map[122];
			agg_result[123] <= discount_cl[123] * bit_map[123];
			agg_result[124] <= discount_cl[124] * bit_map[124];
			agg_result[125] <= discount_cl[125] * bit_map[125];
			agg_result[126] <= discount_cl[126] * bit_map[126];
			agg_result[127] <= discount_cl[127] * bit_map[127];
			agg_result[128] <= discount_cl[128] * bit_map[128];
			agg_result[129] <= discount_cl[129] * bit_map[129];
			agg_result[130] <= discount_cl[130] * bit_map[130];
			agg_result[131] <= discount_cl[131] * bit_map[131];
			agg_result[132] <= discount_cl[132] * bit_map[132];
			agg_result[133] <= discount_cl[133] * bit_map[133];
			agg_result[134] <= discount_cl[134] * bit_map[134];
			agg_result[135] <= discount_cl[135] * bit_map[135];
			agg_result[136] <= discount_cl[136] * bit_map[136];
			agg_result[137] <= discount_cl[137] * bit_map[137];
			agg_result[138] <= discount_cl[138] * bit_map[138];
			agg_result[139] <= discount_cl[139] * bit_map[139];
			agg_result[140] <= discount_cl[140] * bit_map[140];
			agg_result[141] <= discount_cl[141] * bit_map[141];
			agg_result[142] <= discount_cl[142] * bit_map[142];
			agg_result[143] <= discount_cl[143] * bit_map[143];
			agg_result[144] <= discount_cl[144] * bit_map[144];
			agg_result[145] <= discount_cl[145] * bit_map[145];
			agg_result[146] <= discount_cl[146] * bit_map[146];
			agg_result[147] <= discount_cl[147] * bit_map[147];
			agg_result[148] <= discount_cl[148] * bit_map[148];
			agg_result[149] <= discount_cl[149] * bit_map[149];
			agg_result[150] <= discount_cl[150] * bit_map[150];
			agg_result[151] <= discount_cl[151] * bit_map[151];
			agg_result[152] <= discount_cl[152] * bit_map[152];
			agg_result[153] <= discount_cl[153] * bit_map[153];
			agg_result[154] <= discount_cl[154] * bit_map[154];
			agg_result[155] <= discount_cl[155] * bit_map[155];
			agg_result[156] <= discount_cl[156] * bit_map[156];
			agg_result[157] <= discount_cl[157] * bit_map[157];
			agg_result[158] <= discount_cl[158] * bit_map[158];
			agg_result[159] <= discount_cl[159] * bit_map[159];
			agg_result[160] <= discount_cl[160] * bit_map[160];
			agg_result[161] <= discount_cl[161] * bit_map[161];
			agg_result[162] <= discount_cl[162] * bit_map[162];
			agg_result[163] <= discount_cl[163] * bit_map[163];
			agg_result[164] <= discount_cl[164] * bit_map[164];
			agg_result[165] <= discount_cl[165] * bit_map[165];
			agg_result[166] <= discount_cl[166] * bit_map[166];
			agg_result[167] <= discount_cl[167] * bit_map[167];
			agg_result[168] <= discount_cl[168] * bit_map[168];
			agg_result[169] <= discount_cl[169] * bit_map[169];
			agg_result[170] <= discount_cl[170] * bit_map[170];
			agg_result[171] <= discount_cl[171] * bit_map[171];
			agg_result[172] <= discount_cl[172] * bit_map[172];
			agg_result[173] <= discount_cl[173] * bit_map[173];
			agg_result[174] <= discount_cl[174] * bit_map[174];
			agg_result[175] <= discount_cl[175] * bit_map[175];
			agg_result[176] <= discount_cl[176] * bit_map[176];
			agg_result[177] <= discount_cl[177] * bit_map[177];
			agg_result[178] <= discount_cl[178] * bit_map[178];
			agg_result[179] <= discount_cl[179] * bit_map[179];
			agg_result[180] <= discount_cl[180] * bit_map[180];
			agg_result[181] <= discount_cl[181] * bit_map[181];
			agg_result[182] <= discount_cl[182] * bit_map[182];
			agg_result[183] <= discount_cl[183] * bit_map[183];
			agg_result[184] <= discount_cl[184] * bit_map[184];
			agg_result[185] <= discount_cl[185] * bit_map[185];
			agg_result[186] <= discount_cl[186] * bit_map[186];
			agg_result[187] <= discount_cl[187] * bit_map[187];
			agg_result[188] <= discount_cl[188] * bit_map[188];
			agg_result[189] <= discount_cl[189] * bit_map[189];
			agg_result[190] <= discount_cl[190] * bit_map[190];
			agg_result[191] <= discount_cl[191] * bit_map[191];
			agg_result[192] <= discount_cl[192] * bit_map[192];
			agg_result[193] <= discount_cl[193] * bit_map[193];
			agg_result[194] <= discount_cl[194] * bit_map[194];
			agg_result[195] <= discount_cl[195] * bit_map[195];
			agg_result[196] <= discount_cl[196] * bit_map[196];
			agg_result[197] <= discount_cl[197] * bit_map[197];
			agg_result[198] <= discount_cl[198] * bit_map[198];
			agg_result[199] <= discount_cl[199] * bit_map[199];
			agg_result[200] <= discount_cl[200] * bit_map[200];
			agg_result[201] <= discount_cl[201] * bit_map[201];
			agg_result[202] <= discount_cl[202] * bit_map[202];
			agg_result[203] <= discount_cl[203] * bit_map[203];
			agg_result[204] <= discount_cl[204] * bit_map[204];
			agg_result[205] <= discount_cl[205] * bit_map[205];
			agg_result[206] <= discount_cl[206] * bit_map[206];
			agg_result[207] <= discount_cl[207] * bit_map[207];
			agg_result[208] <= discount_cl[208] * bit_map[208];
			agg_result[209] <= discount_cl[209] * bit_map[209];
			agg_result[210] <= discount_cl[210] * bit_map[210];
			agg_result[211] <= discount_cl[211] * bit_map[211];
			agg_result[212] <= discount_cl[212] * bit_map[212];
			agg_result[213] <= discount_cl[213] * bit_map[213];
			agg_result[214] <= discount_cl[214] * bit_map[214];
			agg_result[215] <= discount_cl[215] * bit_map[215];
			agg_result[216] <= discount_cl[216] * bit_map[216];
			agg_result[217] <= discount_cl[217] * bit_map[217];
			agg_result[218] <= discount_cl[218] * bit_map[218];
			agg_result[219] <= discount_cl[219] * bit_map[219];
			agg_result[220] <= discount_cl[220] * bit_map[220];
			agg_result[221] <= discount_cl[221] * bit_map[221];
			agg_result[222] <= discount_cl[222] * bit_map[222];
			agg_result[223] <= discount_cl[223] * bit_map[223];
			agg_result[224] <= discount_cl[224] * bit_map[224];
			agg_result[225] <= discount_cl[225] * bit_map[225];
			agg_result[226] <= discount_cl[226] * bit_map[226];
			agg_result[227] <= discount_cl[227] * bit_map[227];
			agg_result[228] <= discount_cl[228] * bit_map[228];
			agg_result[229] <= discount_cl[229] * bit_map[229];
			agg_result[230] <= discount_cl[230] * bit_map[230];
			agg_result[231] <= discount_cl[231] * bit_map[231];
			agg_result[232] <= discount_cl[232] * bit_map[232];
			agg_result[233] <= discount_cl[233] * bit_map[233];
			agg_result[234] <= discount_cl[234] * bit_map[234];
			agg_result[235] <= discount_cl[235] * bit_map[235];
			agg_result[236] <= discount_cl[236] * bit_map[236];
			agg_result[237] <= discount_cl[237] * bit_map[237];
			agg_result[238] <= discount_cl[238] * bit_map[238];
			agg_result[239] <= discount_cl[239] * bit_map[239];
			agg_result[240] <= discount_cl[240] * bit_map[240];
			agg_result[241] <= discount_cl[241] * bit_map[241];
			agg_result[242] <= discount_cl[242] * bit_map[242];
			agg_result[243] <= discount_cl[243] * bit_map[243];
			agg_result[244] <= discount_cl[244] * bit_map[244];
			agg_result[245] <= discount_cl[245] * bit_map[245];
			agg_result[246] <= discount_cl[246] * bit_map[246];
			agg_result[247] <= discount_cl[247] * bit_map[247];
			agg_result[248] <= discount_cl[248] * bit_map[248];
			agg_result[249] <= discount_cl[249] * bit_map[249];
			agg_result[250] <= discount_cl[250] * bit_map[250];
			agg_result[251] <= discount_cl[251] * bit_map[251];
			agg_result[252] <= discount_cl[252] * bit_map[252];
			agg_result[253] <= discount_cl[253] * bit_map[253];
			agg_result[254] <= discount_cl[254] * bit_map[254];
			agg_result[255] <= discount_cl[255] * bit_map[255];
			agg_result[256] <= discount_cl[256] * bit_map[256];
			agg_result[257] <= discount_cl[257] * bit_map[257];
			agg_result[258] <= discount_cl[258] * bit_map[258];
			agg_result[259] <= discount_cl[259] * bit_map[259];
			agg_result[260] <= discount_cl[260] * bit_map[260];
			agg_result[261] <= discount_cl[261] * bit_map[261];
			agg_result[262] <= discount_cl[262] * bit_map[262];
			agg_result[263] <= discount_cl[263] * bit_map[263];
			agg_result[264] <= discount_cl[264] * bit_map[264];
			agg_result[265] <= discount_cl[265] * bit_map[265];
			agg_result[266] <= discount_cl[266] * bit_map[266];
			agg_result[267] <= discount_cl[267] * bit_map[267];
			agg_result[268] <= discount_cl[268] * bit_map[268];
			agg_result[269] <= discount_cl[269] * bit_map[269];
			agg_result[270] <= discount_cl[270] * bit_map[270];
			agg_result[271] <= discount_cl[271] * bit_map[271];
			agg_result[272] <= discount_cl[272] * bit_map[272];
			agg_result[273] <= discount_cl[273] * bit_map[273];
			agg_result[274] <= discount_cl[274] * bit_map[274];
			agg_result[275] <= discount_cl[275] * bit_map[275];
			agg_result[276] <= discount_cl[276] * bit_map[276];
			agg_result[277] <= discount_cl[277] * bit_map[277];
			agg_result[278] <= discount_cl[278] * bit_map[278];
			agg_result[279] <= discount_cl[279] * bit_map[279];
			agg_result[280] <= discount_cl[280] * bit_map[280];
			agg_result[281] <= discount_cl[281] * bit_map[281];
			agg_result[282] <= discount_cl[282] * bit_map[282];
			agg_result[283] <= discount_cl[283] * bit_map[283];
			agg_result[284] <= discount_cl[284] * bit_map[284];
			agg_result[285] <= discount_cl[285] * bit_map[285];
			agg_result[286] <= discount_cl[286] * bit_map[286];
			agg_result[287] <= discount_cl[287] * bit_map[287];
			agg_result[288] <= discount_cl[288] * bit_map[288];
			agg_result[289] <= discount_cl[289] * bit_map[289];
			agg_result[290] <= discount_cl[290] * bit_map[290];
			agg_result[291] <= discount_cl[291] * bit_map[291];
			agg_result[292] <= discount_cl[292] * bit_map[292];
			agg_result[293] <= discount_cl[293] * bit_map[293];
			agg_result[294] <= discount_cl[294] * bit_map[294];
			agg_result[295] <= discount_cl[295] * bit_map[295];
			agg_result[296] <= discount_cl[296] * bit_map[296];
			agg_result[297] <= discount_cl[297] * bit_map[297];
			agg_result[298] <= discount_cl[298] * bit_map[298];
			agg_result[299] <= discount_cl[299] * bit_map[299];
			agg_result[300] <= discount_cl[300] * bit_map[300];
			agg_result[301] <= discount_cl[301] * bit_map[301];
			agg_result[302] <= discount_cl[302] * bit_map[302];
			agg_result[303] <= discount_cl[303] * bit_map[303];
			agg_result[304] <= discount_cl[304] * bit_map[304];
			agg_result[305] <= discount_cl[305] * bit_map[305];
			agg_result[306] <= discount_cl[306] * bit_map[306];
			agg_result[307] <= discount_cl[307] * bit_map[307];
			agg_result[308] <= discount_cl[308] * bit_map[308];
			agg_result[309] <= discount_cl[309] * bit_map[309];
			agg_result[310] <= discount_cl[310] * bit_map[310];
			agg_result[311] <= discount_cl[311] * bit_map[311];
			agg_result[312] <= discount_cl[312] * bit_map[312];
			agg_result[313] <= discount_cl[313] * bit_map[313];
			agg_result[314] <= discount_cl[314] * bit_map[314];
			agg_result[315] <= discount_cl[315] * bit_map[315];
			agg_result[316] <= discount_cl[316] * bit_map[316];
			agg_result[317] <= discount_cl[317] * bit_map[317];
			agg_result[318] <= discount_cl[318] * bit_map[318];
			agg_result[319] <= discount_cl[319] * bit_map[319];
			agg_result[320] <= discount_cl[320] * bit_map[320];
			agg_result[321] <= discount_cl[321] * bit_map[321];
			agg_result[322] <= discount_cl[322] * bit_map[322];
			agg_result[323] <= discount_cl[323] * bit_map[323];
			agg_result[324] <= discount_cl[324] * bit_map[324];
			agg_result[325] <= discount_cl[325] * bit_map[325];
			agg_result[326] <= discount_cl[326] * bit_map[326];
			agg_result[327] <= discount_cl[327] * bit_map[327];
			agg_result[328] <= discount_cl[328] * bit_map[328];
			agg_result[329] <= discount_cl[329] * bit_map[329];
			agg_result[330] <= discount_cl[330] * bit_map[330];
			agg_result[331] <= discount_cl[331] * bit_map[331];
			agg_result[332] <= discount_cl[332] * bit_map[332];
			agg_result[333] <= discount_cl[333] * bit_map[333];
			agg_result[334] <= discount_cl[334] * bit_map[334];
			agg_result[335] <= discount_cl[335] * bit_map[335];
			agg_result[336] <= discount_cl[336] * bit_map[336];
			agg_result[337] <= discount_cl[337] * bit_map[337];
			agg_result[338] <= discount_cl[338] * bit_map[338];
			agg_result[339] <= discount_cl[339] * bit_map[339];
			agg_result[340] <= discount_cl[340] * bit_map[340];
			agg_result[341] <= discount_cl[341] * bit_map[341];
			agg_result[342] <= discount_cl[342] * bit_map[342];
			agg_result[343] <= discount_cl[343] * bit_map[343];
			agg_result[344] <= discount_cl[344] * bit_map[344];
			agg_result[345] <= discount_cl[345] * bit_map[345];
			agg_result[346] <= discount_cl[346] * bit_map[346];
			agg_result[347] <= discount_cl[347] * bit_map[347];
			agg_result[348] <= discount_cl[348] * bit_map[348];
			agg_result[349] <= discount_cl[349] * bit_map[349];
			agg_result[350] <= discount_cl[350] * bit_map[350];
			agg_result[351] <= discount_cl[351] * bit_map[351];
			agg_result[352] <= discount_cl[352] * bit_map[352];
			agg_result[353] <= discount_cl[353] * bit_map[353];
			agg_result[354] <= discount_cl[354] * bit_map[354];
			agg_result[355] <= discount_cl[355] * bit_map[355];
			agg_result[356] <= discount_cl[356] * bit_map[356];
			agg_result[357] <= discount_cl[357] * bit_map[357];
			agg_result[358] <= discount_cl[358] * bit_map[358];
			agg_result[359] <= discount_cl[359] * bit_map[359];
			agg_result[360] <= discount_cl[360] * bit_map[360];
			agg_result[361] <= discount_cl[361] * bit_map[361];
			agg_result[362] <= discount_cl[362] * bit_map[362];
			agg_result[363] <= discount_cl[363] * bit_map[363];
			agg_result[364] <= discount_cl[364] * bit_map[364];
			agg_result[365] <= discount_cl[365] * bit_map[365];
			agg_result[366] <= discount_cl[366] * bit_map[366];
			agg_result[367] <= discount_cl[367] * bit_map[367];
			agg_result[368] <= discount_cl[368] * bit_map[368];
			agg_result[369] <= discount_cl[369] * bit_map[369];
			agg_result[370] <= discount_cl[370] * bit_map[370];
			agg_result[371] <= discount_cl[371] * bit_map[371];
			agg_result[372] <= discount_cl[372] * bit_map[372];
			agg_result[373] <= discount_cl[373] * bit_map[373];
			agg_result[374] <= discount_cl[374] * bit_map[374];
			agg_result[375] <= discount_cl[375] * bit_map[375];
			agg_result[376] <= discount_cl[376] * bit_map[376];
			agg_result[377] <= discount_cl[377] * bit_map[377];
			agg_result[378] <= discount_cl[378] * bit_map[378];
			agg_result[379] <= discount_cl[379] * bit_map[379];
			agg_result[380] <= discount_cl[380] * bit_map[380];
			agg_result[381] <= discount_cl[381] * bit_map[381];
			agg_result[382] <= discount_cl[382] * bit_map[382];
			agg_result[383] <= discount_cl[383] * bit_map[383];
			agg_result[384] <= discount_cl[384] * bit_map[384];
			agg_result[385] <= discount_cl[385] * bit_map[385];
			agg_result[386] <= discount_cl[386] * bit_map[386];
			agg_result[387] <= discount_cl[387] * bit_map[387];
			agg_result[388] <= discount_cl[388] * bit_map[388];
			agg_result[389] <= discount_cl[389] * bit_map[389];
			agg_result[390] <= discount_cl[390] * bit_map[390];
			agg_result[391] <= discount_cl[391] * bit_map[391];
			agg_result[392] <= discount_cl[392] * bit_map[392];
			agg_result[393] <= discount_cl[393] * bit_map[393];
			agg_result[394] <= discount_cl[394] * bit_map[394];
			agg_result[395] <= discount_cl[395] * bit_map[395];
			agg_result[396] <= discount_cl[396] * bit_map[396];
			agg_result[397] <= discount_cl[397] * bit_map[397];
			agg_result[398] <= discount_cl[398] * bit_map[398];
			agg_result[399] <= discount_cl[399] * bit_map[399];
			agg_result[400] <= discount_cl[400] * bit_map[400];
			agg_result[401] <= discount_cl[401] * bit_map[401];
			agg_result[402] <= discount_cl[402] * bit_map[402];
			agg_result[403] <= discount_cl[403] * bit_map[403];
			agg_result[404] <= discount_cl[404] * bit_map[404];
			agg_result[405] <= discount_cl[405] * bit_map[405];
			agg_result[406] <= discount_cl[406] * bit_map[406];
			agg_result[407] <= discount_cl[407] * bit_map[407];
			agg_result[408] <= discount_cl[408] * bit_map[408];
			agg_result[409] <= discount_cl[409] * bit_map[409];
			agg_result[410] <= discount_cl[410] * bit_map[410];
			agg_result[411] <= discount_cl[411] * bit_map[411];
			agg_result[412] <= discount_cl[412] * bit_map[412];
			agg_result[413] <= discount_cl[413] * bit_map[413];
			agg_result[414] <= discount_cl[414] * bit_map[414];
			agg_result[415] <= discount_cl[415] * bit_map[415];
			agg_result[416] <= discount_cl[416] * bit_map[416];
			agg_result[417] <= discount_cl[417] * bit_map[417];
			agg_result[418] <= discount_cl[418] * bit_map[418];
			agg_result[419] <= discount_cl[419] * bit_map[419];
			agg_result[420] <= discount_cl[420] * bit_map[420];
			agg_result[421] <= discount_cl[421] * bit_map[421];
			agg_result[422] <= discount_cl[422] * bit_map[422];
			agg_result[423] <= discount_cl[423] * bit_map[423];
			agg_result[424] <= discount_cl[424] * bit_map[424];
			agg_result[425] <= discount_cl[425] * bit_map[425];
			agg_result[426] <= discount_cl[426] * bit_map[426];
			agg_result[427] <= discount_cl[427] * bit_map[427];
			agg_result[428] <= discount_cl[428] * bit_map[428];
			agg_result[429] <= discount_cl[429] * bit_map[429];
			agg_result[430] <= discount_cl[430] * bit_map[430];
			agg_result[431] <= discount_cl[431] * bit_map[431];
			agg_result[432] <= discount_cl[432] * bit_map[432];
			agg_result[433] <= discount_cl[433] * bit_map[433];
			agg_result[434] <= discount_cl[434] * bit_map[434];
			agg_result[435] <= discount_cl[435] * bit_map[435];
			agg_result[436] <= discount_cl[436] * bit_map[436];
			agg_result[437] <= discount_cl[437] * bit_map[437];
			agg_result[438] <= discount_cl[438] * bit_map[438];
			agg_result[439] <= discount_cl[439] * bit_map[439];
			agg_result[440] <= discount_cl[440] * bit_map[440];
			agg_result[441] <= discount_cl[441] * bit_map[441];
			agg_result[442] <= discount_cl[442] * bit_map[442];
			agg_result[443] <= discount_cl[443] * bit_map[443];
			agg_result[444] <= discount_cl[444] * bit_map[444];
			agg_result[445] <= discount_cl[445] * bit_map[445];
			agg_result[446] <= discount_cl[446] * bit_map[446];
			agg_result[447] <= discount_cl[447] * bit_map[447];
			agg_result[448] <= discount_cl[448] * bit_map[448];
			agg_result[449] <= discount_cl[449] * bit_map[449];
			agg_result[450] <= discount_cl[450] * bit_map[450];
			agg_result[451] <= discount_cl[451] * bit_map[451];
			agg_result[452] <= discount_cl[452] * bit_map[452];
			agg_result[453] <= discount_cl[453] * bit_map[453];
			agg_result[454] <= discount_cl[454] * bit_map[454];
			agg_result[455] <= discount_cl[455] * bit_map[455];
			agg_result[456] <= discount_cl[456] * bit_map[456];
			agg_result[457] <= discount_cl[457] * bit_map[457];
			agg_result[458] <= discount_cl[458] * bit_map[458];
			agg_result[459] <= discount_cl[459] * bit_map[459];
			agg_result[460] <= discount_cl[460] * bit_map[460];
			agg_result[461] <= discount_cl[461] * bit_map[461];
			agg_result[462] <= discount_cl[462] * bit_map[462];
			agg_result[463] <= discount_cl[463] * bit_map[463];
			agg_result[464] <= discount_cl[464] * bit_map[464];
			agg_result[465] <= discount_cl[465] * bit_map[465];
			agg_result[466] <= discount_cl[466] * bit_map[466];
			agg_result[467] <= discount_cl[467] * bit_map[467];
			agg_result[468] <= discount_cl[468] * bit_map[468];
			agg_result[469] <= discount_cl[469] * bit_map[469];
			agg_result[470] <= discount_cl[470] * bit_map[470];
			agg_result[471] <= discount_cl[471] * bit_map[471];
			agg_result[472] <= discount_cl[472] * bit_map[472];
			agg_result[473] <= discount_cl[473] * bit_map[473];
			agg_result[474] <= discount_cl[474] * bit_map[474];
			agg_result[475] <= discount_cl[475] * bit_map[475];
			agg_result[476] <= discount_cl[476] * bit_map[476];
			agg_result[477] <= discount_cl[477] * bit_map[477];
			agg_result[478] <= discount_cl[478] * bit_map[478];
			agg_result[479] <= discount_cl[479] * bit_map[479];
			agg_result[480] <= discount_cl[480] * bit_map[480];
			agg_result[481] <= discount_cl[481] * bit_map[481];
			agg_result[482] <= discount_cl[482] * bit_map[482];
			agg_result[483] <= discount_cl[483] * bit_map[483];
			agg_result[484] <= discount_cl[484] * bit_map[484];
			agg_result[485] <= discount_cl[485] * bit_map[485];
			agg_result[486] <= discount_cl[486] * bit_map[486];
			agg_result[487] <= discount_cl[487] * bit_map[487];
			agg_result[488] <= discount_cl[488] * bit_map[488];
			agg_result[489] <= discount_cl[489] * bit_map[489];
			agg_result[490] <= discount_cl[490] * bit_map[490];
			agg_result[491] <= discount_cl[491] * bit_map[491];
			agg_result[492] <= discount_cl[492] * bit_map[492];
			agg_result[493] <= discount_cl[493] * bit_map[493];
			agg_result[494] <= discount_cl[494] * bit_map[494];
			agg_result[495] <= discount_cl[495] * bit_map[495];
			agg_result[496] <= discount_cl[496] * bit_map[496];
			agg_result[497] <= discount_cl[497] * bit_map[497];
			agg_result[498] <= discount_cl[498] * bit_map[498];
			agg_result[499] <= discount_cl[499] * bit_map[499];
			agg_result[500] <= discount_cl[500] * bit_map[500];
			agg_result[501] <= discount_cl[501] * bit_map[501];
			agg_result[502] <= discount_cl[502] * bit_map[502];
			agg_result[503] <= discount_cl[503] * bit_map[503];
			agg_result[504] <= discount_cl[504] * bit_map[504];
			agg_result[505] <= discount_cl[505] * bit_map[505];
			agg_result[506] <= discount_cl[506] * bit_map[506];
			agg_result[507] <= discount_cl[507] * bit_map[507];
			agg_result[508] <= discount_cl[508] * bit_map[508];
			agg_result[509] <= discount_cl[509] * bit_map[509];
			agg_result[510] <= discount_cl[510] * bit_map[510];
			agg_result[511] <= discount_cl[511] * bit_map[511];									
			processing_done <= 1'b1;
		end	
	end				
endmodule
