//
// Application configuration.
//

// This application doesn't use MPF
//`define MPF_DISABLED 1
`define MPF_CONF_ENABLE_VTP 1

//`define MPF_CONF_VTP_PT_MODE_SOFTWARE_SERVICE
