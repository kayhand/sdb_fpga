`define MPF_CONF_ENABLE_VTP 1